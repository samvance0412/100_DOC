# 100_DOC
100 Days of Code - Log

### Day 1: April 9, 2018 

**Today's Progress**: Started FreeCodeCamp HTML & CSS Challenges, Second set of Data Science coursework, Joined BSIC Impact Incubator Challenge team and read a lot about the different coding languages 

**Thoughts:** Basic concepts are digestible but the definitions can trip me up - difference between Class and style etc. 

### Day 2: April 10, 2018 

**Today's Progress**:

**Thoughts:**
